module MULTI_BIT_NOT_GATE (
	input  a[31:0],
	output b[31:0]);

	not(b[0], a[0]);
	
endmodule
